use ieee.e
